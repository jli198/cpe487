-- intermediate signal declaration
signal p1_out,p2_out,p3_out : std_logic;