entity my_entity is
port(
	port_name_1 : in std_logic;
	port_name_2 : out std_logic;
	port_name_3 : inout std_logic); --do not forget semicolon
end my_entity; -- do not forget this semicolon either