-- for loop
my_label: for index in a_range loop
	sequential stateemnts...
end loop my_label;

-- while loop
my_label: while (condition) loop
	sequential statements...
end loop my_label;