if x = '0' and y = '0' or z = '1' then
	blah; -- some useful statement
	blah; -- some useful statement
end if;
if ( ((x = '0') and (y = '0')) or (z = '1') ) then
	blah; -- some useful statement
	blah; -- some useful statement
end if;