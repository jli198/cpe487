signal mode: bit;
mode<='0','1' after 10ns,'0' after 30ns,'1' after 40ns,'0' after 70ns;